/*
 * Copyright (c) 2024 Eric Fogleman
 * SPDX-License-Identifier: Apache-2.0
 *
 * TT project wrapper for ef_smsdac
 * 1-10 MHz Segmented mismatch-shaping DAC 
 * Input clock at 1-50 MHz 
 * 8-b unsigned input data on ui_in[7:0]; sync'd to clk (oversampled)
 * uo_out[7:0] connect to {8x, 4x, 2x, 1x} weight 3-level DACs
 * uio currently unused (create SPI data interface in future)
 */

`default_nettype none

module tt_um_ejfogleman_smsdac (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
    );

  // uio currently unused.
  assign uio_out = 0;
  assign uio_oe  = 0;

  u_dac_top ef_smsdac_top( 
    .clk(clk), 
    .rst_b(rst_n), 
    .d_in(ui_in[7:0]), 
    .d_out_3(uo_out[7:6]), 
    .d_out_2(uo_out[5:4]), 
    .d_out_1(uo_out[3:2]), 
    .d_out_0(uo_out[1:0]) );

endmodule
